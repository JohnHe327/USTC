
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h0584d263;
    ram_cell[       1] = 32'h0;  // 32'h16b6a656;
    ram_cell[       2] = 32'h0;  // 32'h59eea795;
    ram_cell[       3] = 32'h0;  // 32'h614a26a7;
    ram_cell[       4] = 32'h0;  // 32'hf76711f7;
    ram_cell[       5] = 32'h0;  // 32'h27d5a98a;
    ram_cell[       6] = 32'h0;  // 32'hd15c1026;
    ram_cell[       7] = 32'h0;  // 32'h1adc0762;
    ram_cell[       8] = 32'h0;  // 32'h02d028ba;
    ram_cell[       9] = 32'h0;  // 32'h50525809;
    ram_cell[      10] = 32'h0;  // 32'hc01d2458;
    ram_cell[      11] = 32'h0;  // 32'ha90a9ee6;
    ram_cell[      12] = 32'h0;  // 32'hb41fdf9c;
    ram_cell[      13] = 32'h0;  // 32'h6226ae7a;
    ram_cell[      14] = 32'h0;  // 32'h8d81421a;
    ram_cell[      15] = 32'h0;  // 32'hc33447d1;
    ram_cell[      16] = 32'h0;  // 32'hf384fad4;
    ram_cell[      17] = 32'h0;  // 32'hc5a1f423;
    ram_cell[      18] = 32'h0;  // 32'h4d06c0fe;
    ram_cell[      19] = 32'h0;  // 32'h094750c9;
    ram_cell[      20] = 32'h0;  // 32'hdd6284ba;
    ram_cell[      21] = 32'h0;  // 32'h6c18ad4d;
    ram_cell[      22] = 32'h0;  // 32'h2521587c;
    ram_cell[      23] = 32'h0;  // 32'hbd719deb;
    ram_cell[      24] = 32'h0;  // 32'h36228092;
    ram_cell[      25] = 32'h0;  // 32'h2d59623d;
    ram_cell[      26] = 32'h0;  // 32'h6cb9b4df;
    ram_cell[      27] = 32'h0;  // 32'hc183cc35;
    ram_cell[      28] = 32'h0;  // 32'hb5c24f18;
    ram_cell[      29] = 32'h0;  // 32'h3b548796;
    ram_cell[      30] = 32'h0;  // 32'hfa0181fd;
    ram_cell[      31] = 32'h0;  // 32'h48bba850;
    ram_cell[      32] = 32'h0;  // 32'h0b598b92;
    ram_cell[      33] = 32'h0;  // 32'h9c740718;
    ram_cell[      34] = 32'h0;  // 32'hd46f30ac;
    ram_cell[      35] = 32'h0;  // 32'h17dd92fa;
    ram_cell[      36] = 32'h0;  // 32'ha8492261;
    ram_cell[      37] = 32'h0;  // 32'h16e7e052;
    ram_cell[      38] = 32'h0;  // 32'h5f736768;
    ram_cell[      39] = 32'h0;  // 32'he76c0895;
    ram_cell[      40] = 32'h0;  // 32'h0da6696d;
    ram_cell[      41] = 32'h0;  // 32'ha5701c50;
    ram_cell[      42] = 32'h0;  // 32'h01076808;
    ram_cell[      43] = 32'h0;  // 32'h210243ae;
    ram_cell[      44] = 32'h0;  // 32'h40bbd3b4;
    ram_cell[      45] = 32'h0;  // 32'h87f92471;
    ram_cell[      46] = 32'h0;  // 32'h48b6b18e;
    ram_cell[      47] = 32'h0;  // 32'h55dcff0f;
    ram_cell[      48] = 32'h0;  // 32'hc80e1748;
    ram_cell[      49] = 32'h0;  // 32'h65c0a88b;
    ram_cell[      50] = 32'h0;  // 32'hd81c0a08;
    ram_cell[      51] = 32'h0;  // 32'hc0db9cd8;
    ram_cell[      52] = 32'h0;  // 32'h07aa996f;
    ram_cell[      53] = 32'h0;  // 32'hf3e43082;
    ram_cell[      54] = 32'h0;  // 32'hb8d2e459;
    ram_cell[      55] = 32'h0;  // 32'hc662dc8b;
    ram_cell[      56] = 32'h0;  // 32'hd59ac380;
    ram_cell[      57] = 32'h0;  // 32'he4ff1f1b;
    ram_cell[      58] = 32'h0;  // 32'h5b79e201;
    ram_cell[      59] = 32'h0;  // 32'h6b8af6de;
    ram_cell[      60] = 32'h0;  // 32'h2ce6808a;
    ram_cell[      61] = 32'h0;  // 32'h14d573a7;
    ram_cell[      62] = 32'h0;  // 32'h77275df4;
    ram_cell[      63] = 32'h0;  // 32'h682fa76e;
    ram_cell[      64] = 32'h0;  // 32'hd0c701dc;
    ram_cell[      65] = 32'h0;  // 32'h4aa01543;
    ram_cell[      66] = 32'h0;  // 32'h3d27ac74;
    ram_cell[      67] = 32'h0;  // 32'h0b804eec;
    ram_cell[      68] = 32'h0;  // 32'hfca3d55c;
    ram_cell[      69] = 32'h0;  // 32'hb2ff050b;
    ram_cell[      70] = 32'h0;  // 32'ha05226e8;
    ram_cell[      71] = 32'h0;  // 32'hf92941e5;
    ram_cell[      72] = 32'h0;  // 32'h336f516c;
    ram_cell[      73] = 32'h0;  // 32'hccb1bdd4;
    ram_cell[      74] = 32'h0;  // 32'h6d12e6b3;
    ram_cell[      75] = 32'h0;  // 32'hf48b5ae9;
    ram_cell[      76] = 32'h0;  // 32'h15ecaa6b;
    ram_cell[      77] = 32'h0;  // 32'h6131ffd6;
    ram_cell[      78] = 32'h0;  // 32'hb53827cc;
    ram_cell[      79] = 32'h0;  // 32'hb21bea70;
    ram_cell[      80] = 32'h0;  // 32'h1683f755;
    ram_cell[      81] = 32'h0;  // 32'hdf0a7ac7;
    ram_cell[      82] = 32'h0;  // 32'hd6d48f50;
    ram_cell[      83] = 32'h0;  // 32'hd05da520;
    ram_cell[      84] = 32'h0;  // 32'h270ce165;
    ram_cell[      85] = 32'h0;  // 32'h9b0e8a5c;
    ram_cell[      86] = 32'h0;  // 32'ha9e5e779;
    ram_cell[      87] = 32'h0;  // 32'h2b283821;
    ram_cell[      88] = 32'h0;  // 32'h9438a943;
    ram_cell[      89] = 32'h0;  // 32'h89e8a274;
    ram_cell[      90] = 32'h0;  // 32'h9f78f1da;
    ram_cell[      91] = 32'h0;  // 32'h1a7e6b24;
    ram_cell[      92] = 32'h0;  // 32'h267eb0a4;
    ram_cell[      93] = 32'h0;  // 32'h22ae72f0;
    ram_cell[      94] = 32'h0;  // 32'h25cf6159;
    ram_cell[      95] = 32'h0;  // 32'hff9dfb94;
    ram_cell[      96] = 32'h0;  // 32'h3907d164;
    ram_cell[      97] = 32'h0;  // 32'h14cabd33;
    ram_cell[      98] = 32'h0;  // 32'h46edfaab;
    ram_cell[      99] = 32'h0;  // 32'h01be3bf7;
    ram_cell[     100] = 32'h0;  // 32'h9042d327;
    ram_cell[     101] = 32'h0;  // 32'h84dc7642;
    ram_cell[     102] = 32'h0;  // 32'h3ed92a13;
    ram_cell[     103] = 32'h0;  // 32'h107268b1;
    ram_cell[     104] = 32'h0;  // 32'h2e5520d3;
    ram_cell[     105] = 32'h0;  // 32'h3177c124;
    ram_cell[     106] = 32'h0;  // 32'h2475a030;
    ram_cell[     107] = 32'h0;  // 32'h3b01aec7;
    ram_cell[     108] = 32'h0;  // 32'h51ea7b0e;
    ram_cell[     109] = 32'h0;  // 32'hb792db4b;
    ram_cell[     110] = 32'h0;  // 32'h95448726;
    ram_cell[     111] = 32'h0;  // 32'hd2754336;
    ram_cell[     112] = 32'h0;  // 32'hffdf7cfa;
    ram_cell[     113] = 32'h0;  // 32'h68dfddd9;
    ram_cell[     114] = 32'h0;  // 32'ha40fb020;
    ram_cell[     115] = 32'h0;  // 32'h37ceef6a;
    ram_cell[     116] = 32'h0;  // 32'hdb3a3b22;
    ram_cell[     117] = 32'h0;  // 32'ha4bc0bc4;
    ram_cell[     118] = 32'h0;  // 32'hc318652a;
    ram_cell[     119] = 32'h0;  // 32'h4089dfbd;
    ram_cell[     120] = 32'h0;  // 32'h00273acd;
    ram_cell[     121] = 32'h0;  // 32'hd8b2d985;
    ram_cell[     122] = 32'h0;  // 32'he36e40c9;
    ram_cell[     123] = 32'h0;  // 32'h232c7907;
    ram_cell[     124] = 32'h0;  // 32'h68085342;
    ram_cell[     125] = 32'h0;  // 32'hd36e64e1;
    ram_cell[     126] = 32'h0;  // 32'h6f0d1871;
    ram_cell[     127] = 32'h0;  // 32'h7a32edaa;
    ram_cell[     128] = 32'h0;  // 32'h169a2879;
    ram_cell[     129] = 32'h0;  // 32'h600a2989;
    ram_cell[     130] = 32'h0;  // 32'h249bd5b5;
    ram_cell[     131] = 32'h0;  // 32'hbe674dde;
    ram_cell[     132] = 32'h0;  // 32'h84f3bb8c;
    ram_cell[     133] = 32'h0;  // 32'h3a13d25d;
    ram_cell[     134] = 32'h0;  // 32'h3ee66d1d;
    ram_cell[     135] = 32'h0;  // 32'h3577ca04;
    ram_cell[     136] = 32'h0;  // 32'h1601b437;
    ram_cell[     137] = 32'h0;  // 32'ha1a873c2;
    ram_cell[     138] = 32'h0;  // 32'h513ed589;
    ram_cell[     139] = 32'h0;  // 32'h0ba9b1c3;
    ram_cell[     140] = 32'h0;  // 32'h8e1faef7;
    ram_cell[     141] = 32'h0;  // 32'h0a992c2c;
    ram_cell[     142] = 32'h0;  // 32'hd9ac9b8e;
    ram_cell[     143] = 32'h0;  // 32'h1e5f97f4;
    ram_cell[     144] = 32'h0;  // 32'h115f4392;
    ram_cell[     145] = 32'h0;  // 32'h7938d459;
    ram_cell[     146] = 32'h0;  // 32'h723767e0;
    ram_cell[     147] = 32'h0;  // 32'hf62dc790;
    ram_cell[     148] = 32'h0;  // 32'hc4e57a59;
    ram_cell[     149] = 32'h0;  // 32'h24170fde;
    ram_cell[     150] = 32'h0;  // 32'hd7b14dd5;
    ram_cell[     151] = 32'h0;  // 32'hc0526003;
    ram_cell[     152] = 32'h0;  // 32'ha1523e79;
    ram_cell[     153] = 32'h0;  // 32'hfaeccf2d;
    ram_cell[     154] = 32'h0;  // 32'ha7025a21;
    ram_cell[     155] = 32'h0;  // 32'h38e81b60;
    ram_cell[     156] = 32'h0;  // 32'h05f32313;
    ram_cell[     157] = 32'h0;  // 32'hdd4476b6;
    ram_cell[     158] = 32'h0;  // 32'he16b07e6;
    ram_cell[     159] = 32'h0;  // 32'hd0a85c2b;
    ram_cell[     160] = 32'h0;  // 32'h770e8109;
    ram_cell[     161] = 32'h0;  // 32'h1e80726c;
    ram_cell[     162] = 32'h0;  // 32'h79125250;
    ram_cell[     163] = 32'h0;  // 32'h7eda5752;
    ram_cell[     164] = 32'h0;  // 32'hb402d016;
    ram_cell[     165] = 32'h0;  // 32'hac9195a1;
    ram_cell[     166] = 32'h0;  // 32'hdf25f3dd;
    ram_cell[     167] = 32'h0;  // 32'hc5809414;
    ram_cell[     168] = 32'h0;  // 32'h809fad33;
    ram_cell[     169] = 32'h0;  // 32'hcdca7baf;
    ram_cell[     170] = 32'h0;  // 32'h88064700;
    ram_cell[     171] = 32'h0;  // 32'he652c80d;
    ram_cell[     172] = 32'h0;  // 32'h63e8d97d;
    ram_cell[     173] = 32'h0;  // 32'hafe6284c;
    ram_cell[     174] = 32'h0;  // 32'hd54b5298;
    ram_cell[     175] = 32'h0;  // 32'h5ed703dd;
    ram_cell[     176] = 32'h0;  // 32'hffaf0f56;
    ram_cell[     177] = 32'h0;  // 32'h5aa1b23e;
    ram_cell[     178] = 32'h0;  // 32'h668749e2;
    ram_cell[     179] = 32'h0;  // 32'h0780ee02;
    ram_cell[     180] = 32'h0;  // 32'h24309562;
    ram_cell[     181] = 32'h0;  // 32'h6c4ef1ec;
    ram_cell[     182] = 32'h0;  // 32'heeb9f36c;
    ram_cell[     183] = 32'h0;  // 32'hb4c73a6a;
    ram_cell[     184] = 32'h0;  // 32'h0a3f90f2;
    ram_cell[     185] = 32'h0;  // 32'h5a8212d2;
    ram_cell[     186] = 32'h0;  // 32'h2141c7e4;
    ram_cell[     187] = 32'h0;  // 32'hd600984d;
    ram_cell[     188] = 32'h0;  // 32'ha5bc77ad;
    ram_cell[     189] = 32'h0;  // 32'head21c56;
    ram_cell[     190] = 32'h0;  // 32'hce1798da;
    ram_cell[     191] = 32'h0;  // 32'h29716ac8;
    ram_cell[     192] = 32'h0;  // 32'he3bb5424;
    ram_cell[     193] = 32'h0;  // 32'h7cb364bc;
    ram_cell[     194] = 32'h0;  // 32'h4db1c2f6;
    ram_cell[     195] = 32'h0;  // 32'h3bdf6dbb;
    ram_cell[     196] = 32'h0;  // 32'h3eda709b;
    ram_cell[     197] = 32'h0;  // 32'h5723f035;
    ram_cell[     198] = 32'h0;  // 32'h928e4c38;
    ram_cell[     199] = 32'h0;  // 32'hfd27da8f;
    ram_cell[     200] = 32'h0;  // 32'h481749d7;
    ram_cell[     201] = 32'h0;  // 32'h3a99e3d0;
    ram_cell[     202] = 32'h0;  // 32'haab96ffd;
    ram_cell[     203] = 32'h0;  // 32'heda79192;
    ram_cell[     204] = 32'h0;  // 32'h11c878fa;
    ram_cell[     205] = 32'h0;  // 32'h9098cdbb;
    ram_cell[     206] = 32'h0;  // 32'h0616672c;
    ram_cell[     207] = 32'h0;  // 32'h71a25923;
    ram_cell[     208] = 32'h0;  // 32'he4d3bf62;
    ram_cell[     209] = 32'h0;  // 32'h95c46c15;
    ram_cell[     210] = 32'h0;  // 32'hfd1e519d;
    ram_cell[     211] = 32'h0;  // 32'heb344ea0;
    ram_cell[     212] = 32'h0;  // 32'hdacbf644;
    ram_cell[     213] = 32'h0;  // 32'h82c84ce9;
    ram_cell[     214] = 32'h0;  // 32'h6905b63a;
    ram_cell[     215] = 32'h0;  // 32'h3c02a7b3;
    ram_cell[     216] = 32'h0;  // 32'hc61eefc8;
    ram_cell[     217] = 32'h0;  // 32'hd9894e7c;
    ram_cell[     218] = 32'h0;  // 32'h3b3bacaa;
    ram_cell[     219] = 32'h0;  // 32'hce397ec2;
    ram_cell[     220] = 32'h0;  // 32'he4f56e29;
    ram_cell[     221] = 32'h0;  // 32'hcb939575;
    ram_cell[     222] = 32'h0;  // 32'h7d9fe754;
    ram_cell[     223] = 32'h0;  // 32'h1e89c3de;
    ram_cell[     224] = 32'h0;  // 32'h9e3842f2;
    ram_cell[     225] = 32'h0;  // 32'hf816b5e3;
    ram_cell[     226] = 32'h0;  // 32'h6cbbdc7b;
    ram_cell[     227] = 32'h0;  // 32'h763ca7b2;
    ram_cell[     228] = 32'h0;  // 32'h626f883f;
    ram_cell[     229] = 32'h0;  // 32'h7f7cad90;
    ram_cell[     230] = 32'h0;  // 32'hb67d2b28;
    ram_cell[     231] = 32'h0;  // 32'hd9515341;
    ram_cell[     232] = 32'h0;  // 32'h145c738f;
    ram_cell[     233] = 32'h0;  // 32'hc37b979e;
    ram_cell[     234] = 32'h0;  // 32'h7ea12c70;
    ram_cell[     235] = 32'h0;  // 32'haa0d7848;
    ram_cell[     236] = 32'h0;  // 32'hf3524861;
    ram_cell[     237] = 32'h0;  // 32'h9786c7f9;
    ram_cell[     238] = 32'h0;  // 32'hd9a6c269;
    ram_cell[     239] = 32'h0;  // 32'h65f906cc;
    ram_cell[     240] = 32'h0;  // 32'hf16b0c2d;
    ram_cell[     241] = 32'h0;  // 32'hbbcdde68;
    ram_cell[     242] = 32'h0;  // 32'h22f1944e;
    ram_cell[     243] = 32'h0;  // 32'hfd50225e;
    ram_cell[     244] = 32'h0;  // 32'hf0a67e0c;
    ram_cell[     245] = 32'h0;  // 32'ha4c1b503;
    ram_cell[     246] = 32'h0;  // 32'h107eed31;
    ram_cell[     247] = 32'h0;  // 32'h830560f1;
    ram_cell[     248] = 32'h0;  // 32'h0c56ead5;
    ram_cell[     249] = 32'h0;  // 32'hc4ce8f5f;
    ram_cell[     250] = 32'h0;  // 32'hd8e65d07;
    ram_cell[     251] = 32'h0;  // 32'h9d28f99b;
    ram_cell[     252] = 32'h0;  // 32'h7242652d;
    ram_cell[     253] = 32'h0;  // 32'h2eab0869;
    ram_cell[     254] = 32'h0;  // 32'hdbadf15e;
    ram_cell[     255] = 32'h0;  // 32'hd2035a3d;
    // src matrix A
    ram_cell[     256] = 32'ha8f441b3;
    ram_cell[     257] = 32'hc9802245;
    ram_cell[     258] = 32'h084f2a75;
    ram_cell[     259] = 32'h89503aa2;
    ram_cell[     260] = 32'hb1af638d;
    ram_cell[     261] = 32'hd60778d0;
    ram_cell[     262] = 32'h2c735a26;
    ram_cell[     263] = 32'h4bc61567;
    ram_cell[     264] = 32'h819a631f;
    ram_cell[     265] = 32'h3458615f;
    ram_cell[     266] = 32'hb6b1bf10;
    ram_cell[     267] = 32'h4c87d578;
    ram_cell[     268] = 32'h9ffbaa3a;
    ram_cell[     269] = 32'h728e5d05;
    ram_cell[     270] = 32'haff48e81;
    ram_cell[     271] = 32'hc4fa5aa0;
    ram_cell[     272] = 32'h1b6adc99;
    ram_cell[     273] = 32'h377bf3af;
    ram_cell[     274] = 32'hbc7fcd8b;
    ram_cell[     275] = 32'hadc8c531;
    ram_cell[     276] = 32'h57b56d31;
    ram_cell[     277] = 32'h0119ab9e;
    ram_cell[     278] = 32'hdccddfa7;
    ram_cell[     279] = 32'hd18b38dc;
    ram_cell[     280] = 32'h4a9accc1;
    ram_cell[     281] = 32'hf0a410b1;
    ram_cell[     282] = 32'heb765db3;
    ram_cell[     283] = 32'h4e353051;
    ram_cell[     284] = 32'h6b787fa2;
    ram_cell[     285] = 32'hd3fce582;
    ram_cell[     286] = 32'h25b5256d;
    ram_cell[     287] = 32'hb13e6633;
    ram_cell[     288] = 32'h6a9a3783;
    ram_cell[     289] = 32'hffe4a2e1;
    ram_cell[     290] = 32'h988388bd;
    ram_cell[     291] = 32'h0500ebdd;
    ram_cell[     292] = 32'h399bb4f9;
    ram_cell[     293] = 32'hffed79f6;
    ram_cell[     294] = 32'ha8ad84c2;
    ram_cell[     295] = 32'h7a4fd6d1;
    ram_cell[     296] = 32'h65b346fb;
    ram_cell[     297] = 32'h574afdf5;
    ram_cell[     298] = 32'h67df28c6;
    ram_cell[     299] = 32'h0b82eaa2;
    ram_cell[     300] = 32'hd2c6be86;
    ram_cell[     301] = 32'hd2a43e11;
    ram_cell[     302] = 32'h5ba4bdf6;
    ram_cell[     303] = 32'h6a5ad18b;
    ram_cell[     304] = 32'h31ee95eb;
    ram_cell[     305] = 32'h1375cd1b;
    ram_cell[     306] = 32'hf6132a24;
    ram_cell[     307] = 32'he47c3d13;
    ram_cell[     308] = 32'h88f03efe;
    ram_cell[     309] = 32'hf024ab9d;
    ram_cell[     310] = 32'hd7763a38;
    ram_cell[     311] = 32'h66fca544;
    ram_cell[     312] = 32'h267b88d7;
    ram_cell[     313] = 32'he7ddb600;
    ram_cell[     314] = 32'h105a3981;
    ram_cell[     315] = 32'h549e7d84;
    ram_cell[     316] = 32'h1cb6f500;
    ram_cell[     317] = 32'h5006ce05;
    ram_cell[     318] = 32'h9cbf0dad;
    ram_cell[     319] = 32'hc8d278d1;
    ram_cell[     320] = 32'h8205c0e0;
    ram_cell[     321] = 32'he9a004b9;
    ram_cell[     322] = 32'ha6a652b2;
    ram_cell[     323] = 32'h1380d732;
    ram_cell[     324] = 32'hde29dad4;
    ram_cell[     325] = 32'h9dca3dd5;
    ram_cell[     326] = 32'h5d784b06;
    ram_cell[     327] = 32'h592b00d3;
    ram_cell[     328] = 32'hb78fc3c7;
    ram_cell[     329] = 32'hdbf4fabb;
    ram_cell[     330] = 32'h79fa449b;
    ram_cell[     331] = 32'h01035359;
    ram_cell[     332] = 32'he67fe41e;
    ram_cell[     333] = 32'h09aa93f5;
    ram_cell[     334] = 32'h1c644566;
    ram_cell[     335] = 32'h9609f860;
    ram_cell[     336] = 32'hfeacf12b;
    ram_cell[     337] = 32'h3203adbf;
    ram_cell[     338] = 32'h581cc148;
    ram_cell[     339] = 32'hfa0e4ae6;
    ram_cell[     340] = 32'ha356111f;
    ram_cell[     341] = 32'h6e8cadc3;
    ram_cell[     342] = 32'h5be66cd0;
    ram_cell[     343] = 32'h9e6aa665;
    ram_cell[     344] = 32'ha634daff;
    ram_cell[     345] = 32'h8f494024;
    ram_cell[     346] = 32'h902ecb64;
    ram_cell[     347] = 32'h68708e40;
    ram_cell[     348] = 32'h5e2715cf;
    ram_cell[     349] = 32'hd70a8c44;
    ram_cell[     350] = 32'h8ae47f89;
    ram_cell[     351] = 32'h49e79cf3;
    ram_cell[     352] = 32'hadbf373e;
    ram_cell[     353] = 32'h6b3fbc79;
    ram_cell[     354] = 32'hddb7a992;
    ram_cell[     355] = 32'h3233f113;
    ram_cell[     356] = 32'he8a9457c;
    ram_cell[     357] = 32'h17dac755;
    ram_cell[     358] = 32'hf2064702;
    ram_cell[     359] = 32'hfd74a1db;
    ram_cell[     360] = 32'h5e97de0c;
    ram_cell[     361] = 32'h44f2330d;
    ram_cell[     362] = 32'h596c4f0b;
    ram_cell[     363] = 32'h009d286d;
    ram_cell[     364] = 32'h61d1143d;
    ram_cell[     365] = 32'h71df8402;
    ram_cell[     366] = 32'hce9ab12a;
    ram_cell[     367] = 32'h1f5dc2e4;
    ram_cell[     368] = 32'haa6c9961;
    ram_cell[     369] = 32'h5107bb71;
    ram_cell[     370] = 32'hf87a0b6d;
    ram_cell[     371] = 32'h533cd711;
    ram_cell[     372] = 32'h130ca73b;
    ram_cell[     373] = 32'hf70378b1;
    ram_cell[     374] = 32'h970e0c00;
    ram_cell[     375] = 32'h3e6321d2;
    ram_cell[     376] = 32'haf3d4481;
    ram_cell[     377] = 32'h091559f7;
    ram_cell[     378] = 32'h6cf7e6cd;
    ram_cell[     379] = 32'h9aaa52d0;
    ram_cell[     380] = 32'h5dd24088;
    ram_cell[     381] = 32'h609ea171;
    ram_cell[     382] = 32'h24bc90ce;
    ram_cell[     383] = 32'h1fa6b0d6;
    ram_cell[     384] = 32'h54cb9669;
    ram_cell[     385] = 32'h46841474;
    ram_cell[     386] = 32'h69aba6ee;
    ram_cell[     387] = 32'hf9d67f24;
    ram_cell[     388] = 32'h5b4f1384;
    ram_cell[     389] = 32'h4be13c8e;
    ram_cell[     390] = 32'hd6c176f0;
    ram_cell[     391] = 32'h7a3f2639;
    ram_cell[     392] = 32'hfa0efc50;
    ram_cell[     393] = 32'h4987e1a6;
    ram_cell[     394] = 32'ha771d783;
    ram_cell[     395] = 32'h07f33125;
    ram_cell[     396] = 32'hc7853f4f;
    ram_cell[     397] = 32'hdae0aa45;
    ram_cell[     398] = 32'h06159d19;
    ram_cell[     399] = 32'h648f81d8;
    ram_cell[     400] = 32'h796933a9;
    ram_cell[     401] = 32'h5d873c3b;
    ram_cell[     402] = 32'h8da66294;
    ram_cell[     403] = 32'hb8d17ea8;
    ram_cell[     404] = 32'he467c014;
    ram_cell[     405] = 32'hddb1fa35;
    ram_cell[     406] = 32'ha1640cf2;
    ram_cell[     407] = 32'h7631c544;
    ram_cell[     408] = 32'h55ef8030;
    ram_cell[     409] = 32'h9ea55f43;
    ram_cell[     410] = 32'hc30870c1;
    ram_cell[     411] = 32'h9d87b640;
    ram_cell[     412] = 32'hc98e7fd5;
    ram_cell[     413] = 32'h2667f7a9;
    ram_cell[     414] = 32'hd3c2db17;
    ram_cell[     415] = 32'h6722e5f1;
    ram_cell[     416] = 32'hba31483e;
    ram_cell[     417] = 32'hc052629f;
    ram_cell[     418] = 32'h480328a5;
    ram_cell[     419] = 32'h5223c1ac;
    ram_cell[     420] = 32'hf0b5b7c8;
    ram_cell[     421] = 32'ha93a2829;
    ram_cell[     422] = 32'hedea63e0;
    ram_cell[     423] = 32'hdfc26095;
    ram_cell[     424] = 32'h8efa7a0f;
    ram_cell[     425] = 32'h2c8abb10;
    ram_cell[     426] = 32'h6e32613b;
    ram_cell[     427] = 32'hc2f24f76;
    ram_cell[     428] = 32'h837c86e2;
    ram_cell[     429] = 32'h6a99e012;
    ram_cell[     430] = 32'hd0b8ea9d;
    ram_cell[     431] = 32'ha711bcc0;
    ram_cell[     432] = 32'he1ae3bf9;
    ram_cell[     433] = 32'h3eb19847;
    ram_cell[     434] = 32'hb0ee1d2d;
    ram_cell[     435] = 32'h3ce56f82;
    ram_cell[     436] = 32'ha363b5bd;
    ram_cell[     437] = 32'he67a52c4;
    ram_cell[     438] = 32'he769e92d;
    ram_cell[     439] = 32'h4b3af6e2;
    ram_cell[     440] = 32'hcf011570;
    ram_cell[     441] = 32'h75233a5c;
    ram_cell[     442] = 32'h8a91d166;
    ram_cell[     443] = 32'hac4a2e56;
    ram_cell[     444] = 32'h75afe986;
    ram_cell[     445] = 32'haf9f299d;
    ram_cell[     446] = 32'hc5f9a43e;
    ram_cell[     447] = 32'hb0605e39;
    ram_cell[     448] = 32'hca3e6bce;
    ram_cell[     449] = 32'h69824430;
    ram_cell[     450] = 32'h5fbf18bf;
    ram_cell[     451] = 32'hd2f2eb9b;
    ram_cell[     452] = 32'h09ae58e4;
    ram_cell[     453] = 32'h01158828;
    ram_cell[     454] = 32'h4b47fcb4;
    ram_cell[     455] = 32'h42d95dcd;
    ram_cell[     456] = 32'hea96945e;
    ram_cell[     457] = 32'hc3b4853f;
    ram_cell[     458] = 32'h5fbdc8cd;
    ram_cell[     459] = 32'h9d9b6d85;
    ram_cell[     460] = 32'h2e1422b3;
    ram_cell[     461] = 32'h790fb1d7;
    ram_cell[     462] = 32'h6c5f74ca;
    ram_cell[     463] = 32'hbd5831d6;
    ram_cell[     464] = 32'hf68ab95e;
    ram_cell[     465] = 32'h5d45f5ba;
    ram_cell[     466] = 32'h243799aa;
    ram_cell[     467] = 32'h49b1031a;
    ram_cell[     468] = 32'h4839eb66;
    ram_cell[     469] = 32'hb292fe0e;
    ram_cell[     470] = 32'h5990582c;
    ram_cell[     471] = 32'h1dd1cfdd;
    ram_cell[     472] = 32'h819c8d5d;
    ram_cell[     473] = 32'hf3643b20;
    ram_cell[     474] = 32'h9949d9d5;
    ram_cell[     475] = 32'h72375b36;
    ram_cell[     476] = 32'he456ad77;
    ram_cell[     477] = 32'h40c0c827;
    ram_cell[     478] = 32'h8de6b5b9;
    ram_cell[     479] = 32'h036b3f5a;
    ram_cell[     480] = 32'h870cda46;
    ram_cell[     481] = 32'h819decfa;
    ram_cell[     482] = 32'hb8949c52;
    ram_cell[     483] = 32'h3b8541b7;
    ram_cell[     484] = 32'h1d5d7b69;
    ram_cell[     485] = 32'hdabaafbe;
    ram_cell[     486] = 32'h83a6860d;
    ram_cell[     487] = 32'hcfa41b48;
    ram_cell[     488] = 32'h5be4040f;
    ram_cell[     489] = 32'ha96d4e04;
    ram_cell[     490] = 32'h91ee844c;
    ram_cell[     491] = 32'hcf96a294;
    ram_cell[     492] = 32'hc243389b;
    ram_cell[     493] = 32'h1cd56887;
    ram_cell[     494] = 32'hdba0ac76;
    ram_cell[     495] = 32'h32d282d4;
    ram_cell[     496] = 32'h481cf831;
    ram_cell[     497] = 32'h1f96fcd4;
    ram_cell[     498] = 32'hc7435809;
    ram_cell[     499] = 32'h9e182fe2;
    ram_cell[     500] = 32'h5aba83f6;
    ram_cell[     501] = 32'h99727862;
    ram_cell[     502] = 32'haacbe09a;
    ram_cell[     503] = 32'hd09c26ab;
    ram_cell[     504] = 32'hba78422d;
    ram_cell[     505] = 32'h56099e31;
    ram_cell[     506] = 32'h7b564f96;
    ram_cell[     507] = 32'h10d9dc26;
    ram_cell[     508] = 32'h30e8f67e;
    ram_cell[     509] = 32'hf83bf00f;
    ram_cell[     510] = 32'h89b8ca74;
    ram_cell[     511] = 32'h1dfbda10;
    // src matrix B
    ram_cell[     512] = 32'heaac4288;
    ram_cell[     513] = 32'h001be1f5;
    ram_cell[     514] = 32'h33d24bd6;
    ram_cell[     515] = 32'h6c4ff2c1;
    ram_cell[     516] = 32'h13ee563d;
    ram_cell[     517] = 32'he3fb75f5;
    ram_cell[     518] = 32'h9500b860;
    ram_cell[     519] = 32'hb481d7ec;
    ram_cell[     520] = 32'h40943474;
    ram_cell[     521] = 32'h726490f2;
    ram_cell[     522] = 32'h49d1058f;
    ram_cell[     523] = 32'h8f8cd33b;
    ram_cell[     524] = 32'he2982cf4;
    ram_cell[     525] = 32'h959a0e1d;
    ram_cell[     526] = 32'hb9843470;
    ram_cell[     527] = 32'h85b81085;
    ram_cell[     528] = 32'hf69fc3a8;
    ram_cell[     529] = 32'hb27b106a;
    ram_cell[     530] = 32'h7570e5ad;
    ram_cell[     531] = 32'h0017a92a;
    ram_cell[     532] = 32'h9ab15322;
    ram_cell[     533] = 32'h3fcf7d32;
    ram_cell[     534] = 32'h2e1a3edf;
    ram_cell[     535] = 32'h7748d5bf;
    ram_cell[     536] = 32'heacc9f2d;
    ram_cell[     537] = 32'h65134cef;
    ram_cell[     538] = 32'h322730e0;
    ram_cell[     539] = 32'he57771ac;
    ram_cell[     540] = 32'had7675ba;
    ram_cell[     541] = 32'h8fa20548;
    ram_cell[     542] = 32'h032c8cf1;
    ram_cell[     543] = 32'h159f9914;
    ram_cell[     544] = 32'h1efbb239;
    ram_cell[     545] = 32'h05491048;
    ram_cell[     546] = 32'hdb00ea37;
    ram_cell[     547] = 32'h1b9aa488;
    ram_cell[     548] = 32'h8cb12448;
    ram_cell[     549] = 32'h6d62968b;
    ram_cell[     550] = 32'h5d524b7c;
    ram_cell[     551] = 32'h978c249f;
    ram_cell[     552] = 32'h4cb8b288;
    ram_cell[     553] = 32'hf4dde0ac;
    ram_cell[     554] = 32'h253f7c33;
    ram_cell[     555] = 32'hc811e7e9;
    ram_cell[     556] = 32'h96102ffb;
    ram_cell[     557] = 32'h9cfe3d68;
    ram_cell[     558] = 32'h880abae6;
    ram_cell[     559] = 32'h6925692e;
    ram_cell[     560] = 32'hda588eb0;
    ram_cell[     561] = 32'h61782353;
    ram_cell[     562] = 32'h34ee5d46;
    ram_cell[     563] = 32'h94cfe9e5;
    ram_cell[     564] = 32'h566cd18e;
    ram_cell[     565] = 32'h00fb2617;
    ram_cell[     566] = 32'hc54ebb61;
    ram_cell[     567] = 32'hcb53324e;
    ram_cell[     568] = 32'h0061b00a;
    ram_cell[     569] = 32'h1c03b42a;
    ram_cell[     570] = 32'h9b4b1101;
    ram_cell[     571] = 32'h2ed5dcf4;
    ram_cell[     572] = 32'h60a92ae3;
    ram_cell[     573] = 32'heccbfc7f;
    ram_cell[     574] = 32'hcc994a73;
    ram_cell[     575] = 32'h1e8d6d5b;
    ram_cell[     576] = 32'h51b226cc;
    ram_cell[     577] = 32'h5f8c70e0;
    ram_cell[     578] = 32'haef3d3ad;
    ram_cell[     579] = 32'h1a33372d;
    ram_cell[     580] = 32'h8f3e3bd6;
    ram_cell[     581] = 32'hf3d995ab;
    ram_cell[     582] = 32'h8c94ea00;
    ram_cell[     583] = 32'he5acee58;
    ram_cell[     584] = 32'hdffab545;
    ram_cell[     585] = 32'h0401c68c;
    ram_cell[     586] = 32'h416986fd;
    ram_cell[     587] = 32'h2489ee7f;
    ram_cell[     588] = 32'h79c3d0fb;
    ram_cell[     589] = 32'h44a23ed9;
    ram_cell[     590] = 32'h9ca8fb3e;
    ram_cell[     591] = 32'h0f11f012;
    ram_cell[     592] = 32'hd9527aaf;
    ram_cell[     593] = 32'haa6b90c4;
    ram_cell[     594] = 32'h6da3fee3;
    ram_cell[     595] = 32'h23002696;
    ram_cell[     596] = 32'h042df1ea;
    ram_cell[     597] = 32'h9e46c1ee;
    ram_cell[     598] = 32'h08aa8e6b;
    ram_cell[     599] = 32'hf03dd7d2;
    ram_cell[     600] = 32'h02b2e2e6;
    ram_cell[     601] = 32'h0065db00;
    ram_cell[     602] = 32'h97d7896a;
    ram_cell[     603] = 32'h741ff7cb;
    ram_cell[     604] = 32'hae785518;
    ram_cell[     605] = 32'h4195978b;
    ram_cell[     606] = 32'hbd698913;
    ram_cell[     607] = 32'h129f0c3b;
    ram_cell[     608] = 32'hf4481e88;
    ram_cell[     609] = 32'h486d64ab;
    ram_cell[     610] = 32'h887e865b;
    ram_cell[     611] = 32'h8e81d172;
    ram_cell[     612] = 32'he5440752;
    ram_cell[     613] = 32'hed8ad79a;
    ram_cell[     614] = 32'hb2db6757;
    ram_cell[     615] = 32'h03a17729;
    ram_cell[     616] = 32'h0b68088b;
    ram_cell[     617] = 32'he4a41a7a;
    ram_cell[     618] = 32'h71bc9848;
    ram_cell[     619] = 32'he5ac8513;
    ram_cell[     620] = 32'h16a69059;
    ram_cell[     621] = 32'hc3070da5;
    ram_cell[     622] = 32'h7873a6c5;
    ram_cell[     623] = 32'h476ebdc0;
    ram_cell[     624] = 32'h9a9b555d;
    ram_cell[     625] = 32'h29b2ea47;
    ram_cell[     626] = 32'hb55d615d;
    ram_cell[     627] = 32'hf7263490;
    ram_cell[     628] = 32'h494a8d19;
    ram_cell[     629] = 32'hf71534fb;
    ram_cell[     630] = 32'hea65e509;
    ram_cell[     631] = 32'hd981347d;
    ram_cell[     632] = 32'hfeb79362;
    ram_cell[     633] = 32'h383b501b;
    ram_cell[     634] = 32'h50e01645;
    ram_cell[     635] = 32'h1967814e;
    ram_cell[     636] = 32'h77fc8f41;
    ram_cell[     637] = 32'hc55061e0;
    ram_cell[     638] = 32'h045adb83;
    ram_cell[     639] = 32'h01277952;
    ram_cell[     640] = 32'hd3188c41;
    ram_cell[     641] = 32'hd0e8914e;
    ram_cell[     642] = 32'h22bd2f71;
    ram_cell[     643] = 32'h01a423c0;
    ram_cell[     644] = 32'hc837ecb1;
    ram_cell[     645] = 32'h11c72ad5;
    ram_cell[     646] = 32'h4ee97185;
    ram_cell[     647] = 32'h65edce35;
    ram_cell[     648] = 32'hf52829f7;
    ram_cell[     649] = 32'h3e6d7bee;
    ram_cell[     650] = 32'h00e6b207;
    ram_cell[     651] = 32'h656d49cf;
    ram_cell[     652] = 32'h76703fb9;
    ram_cell[     653] = 32'h84fce34c;
    ram_cell[     654] = 32'hd30a0c33;
    ram_cell[     655] = 32'h22a28bc1;
    ram_cell[     656] = 32'h38797ef2;
    ram_cell[     657] = 32'h2f228f47;
    ram_cell[     658] = 32'h48924ccd;
    ram_cell[     659] = 32'hc7be9f29;
    ram_cell[     660] = 32'hf71641cf;
    ram_cell[     661] = 32'hb86f1e35;
    ram_cell[     662] = 32'ha6c85338;
    ram_cell[     663] = 32'hda480282;
    ram_cell[     664] = 32'h14e38dd9;
    ram_cell[     665] = 32'h36fc40b7;
    ram_cell[     666] = 32'h3a01adb7;
    ram_cell[     667] = 32'hf83d5bbf;
    ram_cell[     668] = 32'h4a17b38b;
    ram_cell[     669] = 32'h44df84af;
    ram_cell[     670] = 32'h950f19ca;
    ram_cell[     671] = 32'h0a4a7a17;
    ram_cell[     672] = 32'h6c3d6735;
    ram_cell[     673] = 32'h0e2fd66f;
    ram_cell[     674] = 32'hc826978e;
    ram_cell[     675] = 32'h50d65874;
    ram_cell[     676] = 32'h036f7d45;
    ram_cell[     677] = 32'ha9dc3b0c;
    ram_cell[     678] = 32'hf97b8871;
    ram_cell[     679] = 32'h3fed469e;
    ram_cell[     680] = 32'h74cf9b82;
    ram_cell[     681] = 32'hcbaec2b4;
    ram_cell[     682] = 32'h0feb654b;
    ram_cell[     683] = 32'h05e766c2;
    ram_cell[     684] = 32'h66c4f826;
    ram_cell[     685] = 32'h331cd777;
    ram_cell[     686] = 32'h55eff30f;
    ram_cell[     687] = 32'hcee1b3ad;
    ram_cell[     688] = 32'ha2f06cca;
    ram_cell[     689] = 32'h739cb7fd;
    ram_cell[     690] = 32'h2c27540d;
    ram_cell[     691] = 32'h443ee483;
    ram_cell[     692] = 32'h16a44142;
    ram_cell[     693] = 32'h9c671fd6;
    ram_cell[     694] = 32'hfbadd49a;
    ram_cell[     695] = 32'ha5885686;
    ram_cell[     696] = 32'hbb2ea96a;
    ram_cell[     697] = 32'h30f7b948;
    ram_cell[     698] = 32'h4dd3b1a1;
    ram_cell[     699] = 32'h99eeb1cf;
    ram_cell[     700] = 32'h76a406d9;
    ram_cell[     701] = 32'hcdaa9cd6;
    ram_cell[     702] = 32'h612b4901;
    ram_cell[     703] = 32'hec03f3fe;
    ram_cell[     704] = 32'h42502d97;
    ram_cell[     705] = 32'hb877c448;
    ram_cell[     706] = 32'hd9d259e8;
    ram_cell[     707] = 32'h69f57b2a;
    ram_cell[     708] = 32'h462aecdc;
    ram_cell[     709] = 32'heb94430b;
    ram_cell[     710] = 32'hf4db1680;
    ram_cell[     711] = 32'h09543203;
    ram_cell[     712] = 32'h26ea4e85;
    ram_cell[     713] = 32'ha4a0d5d9;
    ram_cell[     714] = 32'hc670db91;
    ram_cell[     715] = 32'h754bb606;
    ram_cell[     716] = 32'h21fe2706;
    ram_cell[     717] = 32'h908df89b;
    ram_cell[     718] = 32'hb4a0bde2;
    ram_cell[     719] = 32'h1449f0a0;
    ram_cell[     720] = 32'hbfd50b5c;
    ram_cell[     721] = 32'hc46b26ed;
    ram_cell[     722] = 32'hbaf17d96;
    ram_cell[     723] = 32'h6788edbc;
    ram_cell[     724] = 32'h402f59a6;
    ram_cell[     725] = 32'h10e024d4;
    ram_cell[     726] = 32'h72789751;
    ram_cell[     727] = 32'h7f77e9c8;
    ram_cell[     728] = 32'h4fb81c83;
    ram_cell[     729] = 32'h1586cb2f;
    ram_cell[     730] = 32'h6ca7829e;
    ram_cell[     731] = 32'h39ad4309;
    ram_cell[     732] = 32'hd7522511;
    ram_cell[     733] = 32'hf140ac75;
    ram_cell[     734] = 32'hc63af548;
    ram_cell[     735] = 32'ha6dec50c;
    ram_cell[     736] = 32'h3c6ab41c;
    ram_cell[     737] = 32'h773c8d7e;
    ram_cell[     738] = 32'he3b4c6a7;
    ram_cell[     739] = 32'hc8a22cca;
    ram_cell[     740] = 32'h2d9b98ef;
    ram_cell[     741] = 32'h130d4012;
    ram_cell[     742] = 32'hbf92d888;
    ram_cell[     743] = 32'hbc3f19d4;
    ram_cell[     744] = 32'haed6f26f;
    ram_cell[     745] = 32'h3d5ab0bb;
    ram_cell[     746] = 32'h1689076a;
    ram_cell[     747] = 32'h34775844;
    ram_cell[     748] = 32'h9bedb430;
    ram_cell[     749] = 32'hc0c8aec6;
    ram_cell[     750] = 32'h45789339;
    ram_cell[     751] = 32'h0d7ffeb0;
    ram_cell[     752] = 32'hcc09391d;
    ram_cell[     753] = 32'h15be73eb;
    ram_cell[     754] = 32'h17aa8a30;
    ram_cell[     755] = 32'h08495350;
    ram_cell[     756] = 32'h757aff95;
    ram_cell[     757] = 32'h70c826b1;
    ram_cell[     758] = 32'h02c5ff31;
    ram_cell[     759] = 32'h88344fb5;
    ram_cell[     760] = 32'h93cfd280;
    ram_cell[     761] = 32'h48796358;
    ram_cell[     762] = 32'hd7c42f5b;
    ram_cell[     763] = 32'h37aaae72;
    ram_cell[     764] = 32'h49219ddd;
    ram_cell[     765] = 32'hd3d0e552;
    ram_cell[     766] = 32'h62b21bc6;
    ram_cell[     767] = 32'h1ad38efb;
end

endmodule

