`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: USTC ESLAB
// Engineer: Huang Yifan (hyf15@mail.ustc.edu.cn)
// 
// Design Name: RV32I Core
// Module Name: Instruction Cache
// Tool Versions: Vivado 2017.4.1
// Description: RV32I Instruction Cache
// 
//////////////////////////////////////////////////////////////////////////////////


//  ����˵��
    //  ͬ����д��Cache��ʵ���п��Խ��䵱��ֻ��Cache
    //  debug�˿�����simulationʱ������дָ����Ժ���
// ����
    // clk               ʱ��
    // write_en          debugдʹ��
    // addr              ����ַ
    // debug_addr        debug��д��ַ
    // debug_input       debugдָ��
// ���
    // data              ����ָ��
    // debug_data        debug����ָ��
// ʵ��Ҫ��  
    // �����޸�

// asm file name: btb.S

module InstructionCache(
    input wire clk,
    input wire write_en,
    input wire [31:2] addr, debug_addr,
    input wire [31:0] debug_input,
    output reg [31:0] data, debug_data
);

    // local variable
    wire addr_valid = (addr[31:14] == 18'h0);
    wire debug_addr_valid = (debug_addr[31:14] == 18'h0);
    wire [11:0] dealt_addr = addr[13:2];
    wire [11:0] dealt_debug_addr = debug_addr[13:2];
    // cache content
    reg [31:0] inst_cache[0:4095];


    initial begin
        data = 32'h0;
        debug_data = 32'h0;
        inst_cache[       0] = 32'h00000293;
        inst_cache[       1] = 32'h00000313;
        inst_cache[       2] = 32'h06500393;
        inst_cache[       3] = 32'h00530333;
        inst_cache[       4] = 32'h00128293;
        inst_cache[       5] = 32'hfe729ce3;
        inst_cache[       6] = 32'h00130313;
end

    always@(posedge clk)
    begin
        data <= addr_valid ? inst_cache[dealt_addr] : 32'h0;
        debug_data <= debug_addr_valid ? inst_cache[dealt_debug_addr] : 32'h0;
        if(write_en & debug_addr_valid) 
            inst_cache[dealt_debug_addr] <= debug_input;
    end

endmodule
